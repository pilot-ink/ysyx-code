module top(
	input clk,rst,
  input a,
  input b,
  output f
);
  assign f = a ^ b;
endmodule





