module top(
    input rst,
    input clk
);
    ysyx_24100027_CPU c1(
        .rst(rst),
        .clk(clk)
    );
endmodule

